module decoder(input logic instr[3:0],
		input logic carry,
		output logic [1:0] src_sel, dst_sel,
		output logic src_sel_en, out_3st_en,
		output logic RAM_b_en, ROM_b_en,
		output logic RAM_RW, RAM_WE);

	always_comb
		begin
			
		end
endmodule
